`timescale 1ns / 1ps

module BUFG (O, I);
   output O;
   input I;
endmodule
